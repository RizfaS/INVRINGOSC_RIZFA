magic
tech sky130A
magscale 1 2
timestamp 1729159655
<< nwell >>
rect -189 -803 814 2080
<< nsubdiff >>
rect -153 2010 -93 2044
rect 718 2010 778 2044
rect -153 1984 -119 2010
rect 744 1984 778 2010
rect -153 -733 -119 -708
rect 744 -733 778 -708
rect -153 -767 -93 -733
rect 718 -767 778 -733
<< nsubdiffcont >>
rect -93 2010 718 2044
rect -153 -708 -119 1984
rect 744 -708 778 1984
rect -93 -767 718 -733
<< poly >>
rect -72 1967 24 1983
rect -72 1933 -56 1967
rect -22 1933 24 1967
rect -72 1917 24 1933
rect -6 1907 24 1917
rect 598 1967 694 1983
rect 598 1933 644 1967
rect 678 1933 694 1967
rect 598 1917 694 1933
rect 598 1912 628 1917
rect -72 1273 24 1289
rect 82 1288 282 1390
rect 598 1290 694 1306
rect -72 1239 -56 1273
rect -22 1239 24 1273
rect -72 1223 24 1239
rect -6 1218 24 1223
rect 598 1256 644 1290
rect 678 1256 694 1290
rect 598 1240 694 1256
rect 598 1218 628 1240
rect 615 1199 628 1202
rect 82 594 540 696
rect -6 56 24 76
rect -72 40 24 56
rect -72 6 -56 40
rect -22 6 24 40
rect -72 -10 24 6
rect 598 67 628 73
rect 598 51 690 67
rect 598 17 640 51
rect 674 17 690 51
rect 340 -100 540 2
rect 598 1 690 17
rect -6 -627 24 -587
rect -67 -648 24 -627
rect -67 -682 -52 -648
rect -18 -682 24 -648
rect -67 -693 24 -682
rect 598 -627 628 -622
rect 598 -648 689 -627
rect 598 -682 640 -648
rect 674 -682 689 -648
rect 598 -693 689 -682
rect -52 -698 -18 -693
rect 640 -698 674 -693
<< polycont >>
rect -56 1933 -22 1967
rect 644 1933 678 1967
rect -56 1239 -22 1273
rect 644 1256 678 1290
rect -56 6 -22 40
rect 640 17 674 51
rect -52 -682 -18 -648
rect 640 -682 674 -648
<< locali >>
rect -153 2010 -93 2044
rect 718 2010 778 2044
rect -153 1984 -119 2010
rect 744 1984 778 2010
rect -72 1933 -56 1967
rect -22 1933 -6 1967
rect 628 1933 644 1967
rect 678 1933 694 1967
rect -52 1888 -18 1933
rect 640 1889 674 1933
rect 552 1439 586 1485
rect 524 1405 586 1439
rect -72 1239 -56 1273
rect -22 1239 -6 1273
rect 628 1256 644 1290
rect 678 1256 694 1290
rect -52 1192 -18 1239
rect 640 1193 675 1256
rect 552 745 586 792
rect 526 711 586 745
rect 36 545 96 579
rect 36 498 70 545
rect -52 40 -18 97
rect 640 51 674 96
rect -72 6 -56 40
rect -22 6 -6 40
rect 624 17 640 51
rect 674 17 690 51
rect 36 -149 97 -115
rect 36 -197 71 -149
rect 37 -208 70 -197
rect -52 -648 -18 -578
rect 640 -648 674 -595
rect -18 -682 -2 -648
rect 624 -682 640 -648
rect -52 -698 -18 -682
rect 640 -698 674 -682
rect -153 -733 -119 -708
rect 744 -733 778 -708
rect -153 -767 -93 -733
rect 718 -767 778 -733
<< viali >>
rect -56 1933 -22 1967
rect 644 1933 678 1967
rect 744 1934 778 1968
rect -56 1239 -22 1273
rect 644 1256 678 1290
rect -56 6 -22 40
rect 640 17 674 51
rect -153 -682 -119 -648
rect -52 -682 -18 -648
rect 640 -682 674 -648
<< metal1 >>
rect 732 1973 790 1974
rect -68 1967 -10 1973
rect -68 1933 -56 1967
rect -22 1933 -10 1967
rect -68 1927 -10 1933
rect 632 1968 790 1973
rect 632 1967 744 1968
rect 632 1933 644 1967
rect 678 1934 744 1967
rect 778 1934 790 1968
rect 678 1933 790 1934
rect 632 1928 790 1933
rect 632 1927 690 1928
rect -63 1874 -10 1927
rect -63 1862 70 1874
rect -74 1486 -64 1862
rect -8 1498 70 1862
rect -8 1486 2 1498
rect 288 1439 335 1886
rect 634 1883 680 1927
rect 552 1498 674 1874
rect 546 1445 592 1491
rect 288 1405 380 1439
rect -68 1273 -10 1279
rect -68 1239 -56 1273
rect -22 1239 -10 1273
rect -68 1233 -10 1239
rect -57 1218 -10 1233
rect -57 1180 -12 1218
rect -52 804 26 1180
rect 82 804 92 1180
rect 30 539 116 585
rect 30 486 76 539
rect -52 110 70 486
rect -52 60 -18 110
rect -58 46 -12 60
rect -68 40 -10 46
rect -68 6 -56 40
rect -22 6 -10 40
rect -68 0 -10 6
rect 30 -155 116 -109
rect 288 -115 335 1405
rect 507 1399 593 1445
rect 632 1290 690 1296
rect 632 1256 644 1290
rect 678 1256 690 1290
rect 632 1250 690 1256
rect 634 1235 680 1250
rect 635 1181 680 1235
rect 640 1180 674 1181
rect 552 804 674 1180
rect 546 751 592 804
rect 505 705 592 751
rect 530 110 540 486
rect 596 110 674 486
rect 640 57 674 110
rect 628 51 686 57
rect 628 17 640 51
rect 674 17 686 51
rect 628 11 686 17
rect 242 -149 335 -115
rect 30 -200 76 -155
rect -52 -584 70 -208
rect -52 -588 -18 -584
rect -52 -596 -12 -588
rect 288 -596 335 -149
rect 552 -584 630 -208
rect 686 -584 696 -208
rect -58 -640 -12 -596
rect -154 -642 -12 -640
rect -165 -648 -12 -642
rect 634 -648 680 -584
rect -165 -682 -153 -648
rect -119 -682 -52 -648
rect -18 -682 -2 -648
rect 624 -682 640 -648
rect 674 -682 680 -648
rect -165 -688 -12 -682
rect 634 -688 680 -682
rect -154 -692 -18 -688
rect -52 -698 -18 -692
rect 640 -698 674 -688
<< via1 >>
rect -64 1486 -8 1862
rect 26 804 82 1180
rect 540 110 596 486
rect 630 -584 686 -208
<< metal2 >>
rect -65 1862 -5 1888
rect -65 1486 -64 1862
rect -8 1486 -5 1862
rect -65 1369 -5 1486
rect -65 1313 -63 1369
rect -7 1313 -5 1369
rect -65 -15 -5 1313
rect 628 1371 688 1380
rect 628 1302 688 1311
rect 26 1180 82 1190
rect 26 668 82 804
rect 26 612 596 668
rect 540 486 596 612
rect 540 100 596 110
rect -65 -84 -5 -75
rect 630 -17 686 1302
rect 630 -208 686 -73
rect 630 -594 686 -584
<< via2 >>
rect -63 1313 -7 1369
rect 628 1311 688 1371
rect -65 -75 -5 -15
rect 630 -73 686 -17
<< metal3 >>
rect -68 1371 -2 1374
rect 623 1371 693 1376
rect -68 1369 628 1371
rect -68 1313 -63 1369
rect -7 1313 628 1369
rect -68 1311 628 1313
rect 688 1311 693 1371
rect -68 1308 -2 1311
rect 623 1306 693 1311
rect -70 -15 0 -10
rect 625 -15 691 -12
rect -70 -75 -65 -15
rect -5 -17 691 -15
rect -5 -73 630 -17
rect 686 -73 691 -17
rect -5 -75 691 -73
rect -70 -80 0 -75
rect 625 -78 691 -75
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729147632
transform 1 0 9 0 1 992
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729147632
transform 1 0 9 0 1 -396
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729147632
transform 1 0 613 0 1 -396
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729147632
transform 1 0 613 0 1 298
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729147632
transform 1 0 9 0 1 298
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729147632
transform 1 0 613 0 1 992
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729147632
transform 1 0 613 0 1 1686
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729147632
transform 1 0 9 0 1 1686
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729147632
transform 1 0 311 0 1 1686
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729147632
transform 1 0 311 0 1 992
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729147632
transform 1 0 311 0 1 298
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729147632
transform 1 0 311 0 1 -396
box -323 -300 323 300
<< labels >>
flabel metal2 -38 1419 -38 1419 0 FreeSans 1600 0 0 0 D5
port 0 nsew
flabel metal1 307 1414 307 1414 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal2 56 643 56 643 0 FreeSans 1600 0 0 0 D1
port 2 nsew
flabel metal1 53 522 53 522 0 FreeSans 1600 0 0 0 D2
port 3 nsew
<< end >>
