magic
tech sky130A
magscale 1 2
timestamp 1729240501
<< nmos >>
rect -407 -100 -247 100
rect -189 -100 -29 100
rect 29 -100 189 100
rect 247 -100 407 100
<< ndiff >>
rect -465 88 -407 100
rect -465 -88 -453 88
rect -419 -88 -407 88
rect -465 -100 -407 -88
rect -247 88 -189 100
rect -247 -88 -235 88
rect -201 -88 -189 88
rect -247 -100 -189 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 189 88 247 100
rect 189 -88 201 88
rect 235 -88 247 88
rect 189 -100 247 -88
rect 407 88 465 100
rect 407 -88 419 88
rect 453 -88 465 88
rect 407 -100 465 -88
<< ndiffc >>
rect -453 -88 -419 88
rect -235 -88 -201 88
rect -17 -88 17 88
rect 201 -88 235 88
rect 419 -88 453 88
<< poly >>
rect -407 172 -247 188
rect -407 138 -391 172
rect -263 138 -247 172
rect -407 100 -247 138
rect -189 172 -29 188
rect -189 138 -173 172
rect -45 138 -29 172
rect -189 100 -29 138
rect 29 172 189 188
rect 29 138 45 172
rect 173 138 189 172
rect 29 100 189 138
rect 247 172 407 188
rect 247 138 263 172
rect 391 138 407 172
rect 247 100 407 138
rect -407 -138 -247 -100
rect -407 -172 -391 -138
rect -263 -172 -247 -138
rect -407 -188 -247 -172
rect -189 -138 -29 -100
rect -189 -172 -173 -138
rect -45 -172 -29 -138
rect -189 -188 -29 -172
rect 29 -138 189 -100
rect 29 -172 45 -138
rect 173 -172 189 -138
rect 29 -188 189 -172
rect 247 -138 407 -100
rect 247 -172 263 -138
rect 391 -172 407 -138
rect 247 -188 407 -172
<< polycont >>
rect -391 138 -263 172
rect -173 138 -45 172
rect 45 138 173 172
rect 263 138 391 172
rect -391 -172 -263 -138
rect -173 -172 -45 -138
rect 45 -172 173 -138
rect 263 -172 391 -138
<< locali >>
rect -407 138 -391 172
rect -263 138 -247 172
rect -189 138 -173 172
rect -45 138 -29 172
rect 29 138 45 172
rect 173 138 189 172
rect 247 138 263 172
rect 391 138 407 172
rect -453 88 -419 104
rect -453 -104 -419 -88
rect -235 88 -201 104
rect -235 -104 -201 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 201 88 235 104
rect 201 -104 235 -88
rect 419 88 453 104
rect 419 -104 453 -88
rect -407 -172 -391 -138
rect -263 -172 -247 -138
rect -189 -172 -173 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 173 -172 189 -138
rect 247 -172 263 -138
rect 391 -172 407 -138
<< viali >>
rect -391 138 -263 172
rect -173 138 -45 172
rect 45 138 173 172
rect 263 138 391 172
rect -453 -88 -419 88
rect -235 -88 -201 88
rect -17 -88 17 88
rect 201 -88 235 88
rect 419 -88 453 88
rect -391 -172 -263 -138
rect -173 -172 -45 -138
rect 45 -172 173 -138
rect 263 -172 391 -138
<< metal1 >>
rect -403 172 -251 178
rect -403 138 -391 172
rect -263 138 -251 172
rect -403 132 -251 138
rect -185 172 -33 178
rect -185 138 -173 172
rect -45 138 -33 172
rect -185 132 -33 138
rect 33 172 185 178
rect 33 138 45 172
rect 173 138 185 172
rect 33 132 185 138
rect 251 172 403 178
rect 251 138 263 172
rect 391 138 403 172
rect 251 132 403 138
rect -459 88 -413 100
rect -459 -88 -453 88
rect -419 -88 -413 88
rect -459 -100 -413 -88
rect -241 88 -195 100
rect -241 -88 -235 88
rect -201 -88 -195 88
rect -241 -100 -195 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 195 88 241 100
rect 195 -88 201 88
rect 235 -88 241 88
rect 195 -100 241 -88
rect 413 88 459 100
rect 413 -88 419 88
rect 453 -88 459 88
rect 413 -100 459 -88
rect -403 -138 -251 -132
rect -403 -172 -391 -138
rect -263 -172 -251 -138
rect -403 -178 -251 -172
rect -185 -138 -33 -132
rect -185 -172 -173 -138
rect -45 -172 -33 -138
rect -185 -178 -33 -172
rect 33 -138 185 -132
rect 33 -172 45 -138
rect 173 -172 185 -138
rect 33 -178 185 -172
rect 251 -138 403 -132
rect 251 -172 263 -138
rect 391 -172 403 -138
rect 251 -178 403 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
